module   inverter (a_i, y_o);         
 input  a_i;
output  y_o;
 	assign  y_o  =  ~ a_i;
endmodule